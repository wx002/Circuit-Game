;
v_1_9 n08 0 12 ; 
r_3_9 n08 0 1 ; 
r_5_9 n08 0 1 ; 
.OP ; 
.END ; 
